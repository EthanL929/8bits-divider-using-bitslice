magic
tech tsmc180
timestamp 1673625385
<< metal1 >>
rect 13414 891 13461 903
rect 13513 891 13626 903
rect 13678 891 13791 903
rect 13876 891 13956 903
rect 13348 858 14055 870
rect 12589 825 13197 837
rect 13315 825 14088 837
rect 12523 792 14253 804
rect 11137 759 11217 771
rect 11566 759 14154 771
rect 14173 759 14418 771
rect 10411 726 14550 738
rect 10345 693 14763 705
rect 9388 660 14385 672
rect 14437 660 14715 672
rect 14751 672 14763 693
rect 14751 660 14880 672
rect 7969 627 8016 639
rect 8299 627 14022 639
rect 14074 627 15012 639
rect 15064 627 15177 639
rect 15229 627 15342 639
rect 7903 594 11184 606
rect 11236 594 13428 606
rect 13480 594 14781 606
rect 14800 594 15441 606
rect 7870 561 13527 573
rect 13546 561 14451 573
rect 14470 561 15507 573
rect 6121 528 7125 540
rect 7144 528 13758 540
rect 13810 528 13824 540
rect 13843 528 15309 540
rect 15361 528 15672 540
rect 6055 495 14649 507
rect 14668 495 15573 507
rect 15592 495 15837 507
rect 5098 462 13593 474
rect 13645 462 13692 474
rect 13711 462 14220 474
rect 14272 462 14847 474
rect 14899 462 15243 474
rect 15262 462 15969 474
rect 5032 429 7059 441
rect 7078 429 11481 441
rect 11500 429 15078 441
rect 15097 429 16101 441
rect 4669 396 16233 408
rect 4636 363 16431 375
rect 4009 330 15639 342
rect 15691 330 16530 342
rect 3646 297 16266 309
rect 16285 297 16629 309
rect 16681 297 16761 309
rect 3613 264 16563 276
rect 16582 264 16827 276
rect 2986 231 8346 243
rect 8365 231 13923 243
rect 13975 231 14319 243
rect 14338 231 14484 243
rect 14503 231 14616 243
rect 14635 231 14913 243
rect 14932 231 15804 243
rect 15856 231 16134 243
rect 16153 231 16860 243
rect 2623 198 15408 210
rect 15460 198 15474 210
rect 15526 198 15540 210
rect 15559 198 16002 210
rect 16021 198 16596 210
rect 16648 198 16794 210
rect 16846 198 16959 210
rect 2590 165 15738 177
rect 15757 165 16299 177
rect 16318 165 16497 177
rect 16549 165 17073 177
rect 2029 132 3033 144
rect 3052 132 4056 144
rect 4075 132 7983 144
rect 8035 132 14286 144
rect 14305 132 15870 144
rect 15889 132 16398 144
rect 16450 132 16893 144
rect 16912 132 17040 144
rect 17028 115 17040 132
rect 0 99 327 111
rect 1963 99 9303 111
rect 9322 99 15936 111
rect 15988 99 16068 111
rect 16120 99 16200 111
rect 16252 99 16365 111
rect 16384 99 16464 111
rect 16516 99 16827 111
rect 16879 99 16926 111
rect 16978 99 16992 111
rect 17061 111 17073 165
rect 17061 99 17124 111
rect 0 66 13989 78
rect 14041 66 14979 78
rect 15031 66 15144 78
rect 15196 66 17223 78
rect 0 33 309 45
rect 297 16 309 33
rect 346 33 13179 45
rect 13167 16 13179 33
rect 13216 33 16743 45
rect 15378 16 15390 33
rect 15708 16 15720 33
rect 16731 16 16743 33
rect 16780 33 17106 45
rect 17094 16 17106 33
rect 17143 33 17370 45
rect 17358 16 17370 33
rect 297 -1667 309 -960
rect 429 -1671 441 -960
rect 17160 -978 17172 -960
rect 627 -990 17172 -978
rect 627 -1007 639 -990
rect 17292 -978 17304 -960
rect 17209 -990 17304 -978
rect 17424 -978 17436 -960
rect 17556 -978 17568 -960
rect 17622 -978 17634 -960
rect 17341 -990 17568 -978
rect 17589 -990 17634 -978
rect 676 -1023 10986 -1011
rect 11038 -1023 17487 -1011
rect 17589 -1011 17601 -990
rect 17523 -1023 17601 -1011
rect 610 -1056 8940 -1044
rect 17523 -1044 17535 -1023
rect 8992 -1056 17535 -1044
rect 561 -1089 657 -1077
rect 561 -1106 573 -1089
rect 709 -1089 822 -1077
rect 874 -1089 12141 -1077
rect 12160 -1089 17322 -1077
rect 660 -1122 9963 -1110
rect 660 -1143 672 -1122
rect 10015 -1122 17190 -1110
rect 528 -1155 672 -1143
rect 528 -1601 540 -1155
rect 742 -1155 1251 -1143
rect 1303 -1155 11019 -1143
rect 660 -1188 5673 -1176
rect 561 -1638 573 -1191
rect 594 -1634 606 -1191
rect 627 -1634 639 -1191
rect 660 -1634 672 -1188
rect 5725 -1188 6696 -1176
rect 6748 -1188 9996 -1176
rect 759 -1221 8973 -1209
rect 693 -1634 705 -1224
rect 726 -1634 738 -1224
rect 759 -1634 771 -1221
rect 792 -1254 7719 -1242
rect 792 -1634 804 -1254
rect 825 -1287 6729 -1275
rect 825 -1634 837 -1287
rect 891 -1320 5706 -1308
rect 858 -1634 870 -1323
rect 891 -1634 903 -1320
rect 924 -1353 1284 -1341
rect 495 -1650 573 -1638
rect 495 -1667 507 -1650
rect 330 -1683 441 -1671
rect 330 -1704 342 -1683
rect 924 -1671 936 -1353
rect 577 -1683 936 -1671
rect 280 -1716 342 -1704
rect 379 -1716 657 -1704
rect 231 -1749 294 -1737
rect 231 -1836 243 -1749
rect 891 -1737 903 -1719
rect 346 -1749 903 -1737
rect 297 -1782 855 -1770
rect 198 -1848 243 -1836
rect 198 -1869 210 -1848
rect 264 -1869 276 -1785
rect 297 -1865 309 -1782
rect 412 -1815 822 -1803
rect 330 -1865 342 -1818
rect 363 -1836 375 -1818
rect 363 -1848 426 -1836
rect 478 -1848 789 -1836
rect 165 -1881 210 -1869
rect 231 -1881 276 -1869
rect 165 -1964 177 -1881
rect 231 -1902 243 -1881
rect 379 -1881 756 -1869
rect 198 -1914 243 -1902
rect 198 -1964 210 -1914
rect 280 -1914 723 -1902
rect 231 -1947 690 -1935
rect 231 -1964 243 -1947
<< m2contact >>
rect 13395 888 13414 907
rect 13461 888 13480 907
rect 13494 888 13513 907
rect 13626 888 13645 907
rect 13659 888 13678 907
rect 13791 888 13810 907
rect 13857 888 13876 907
rect 13956 888 13975 907
rect 13329 855 13348 874
rect 14055 855 14074 874
rect 12570 822 12589 841
rect 13197 822 13216 841
rect 13296 822 13315 841
rect 14088 822 14107 841
rect 12504 789 12523 808
rect 14253 789 14272 808
rect 11118 756 11137 775
rect 11217 756 11236 775
rect 11547 756 11566 775
rect 14154 756 14173 775
rect 14418 756 14437 775
rect 10392 723 10411 742
rect 14550 723 14569 742
rect 10326 690 10345 709
rect 9369 657 9388 676
rect 14385 657 14404 676
rect 14418 657 14437 676
rect 14715 657 14734 676
rect 14880 657 14899 676
rect 7950 624 7969 643
rect 8016 624 8035 643
rect 8280 624 8299 643
rect 14022 624 14041 643
rect 14055 624 14074 643
rect 15012 624 15031 643
rect 15045 624 15064 643
rect 15177 624 15196 643
rect 15210 624 15229 643
rect 15342 624 15361 643
rect 7884 591 7903 610
rect 11184 591 11203 610
rect 11217 591 11236 610
rect 13428 591 13447 610
rect 13461 591 13480 610
rect 14781 591 14800 610
rect 15441 591 15460 610
rect 7851 558 7870 577
rect 13527 558 13546 577
rect 14451 558 14470 577
rect 15507 558 15526 577
rect 6102 525 6121 544
rect 7125 525 7144 544
rect 13758 525 13777 544
rect 13791 525 13810 544
rect 13824 525 13843 544
rect 15309 525 15328 544
rect 15342 525 15361 544
rect 15672 525 15691 544
rect 6036 492 6055 511
rect 14649 492 14668 511
rect 15573 492 15592 511
rect 15837 492 15856 511
rect 5079 459 5098 478
rect 13593 459 13612 478
rect 13626 459 13645 478
rect 13692 459 13711 478
rect 14220 459 14239 478
rect 14253 459 14272 478
rect 14847 459 14866 478
rect 14880 459 14899 478
rect 15243 459 15262 478
rect 15969 459 15988 478
rect 5013 426 5032 445
rect 7059 426 7078 445
rect 11481 426 11500 445
rect 15078 426 15097 445
rect 16101 426 16120 445
rect 4650 393 4669 412
rect 16233 393 16252 412
rect 4617 360 4636 379
rect 16431 360 16450 379
rect 3990 327 4009 346
rect 15639 327 15658 346
rect 15672 327 15691 346
rect 16530 327 16549 346
rect 3627 294 3646 313
rect 16266 294 16285 313
rect 16629 294 16648 313
rect 16662 294 16681 313
rect 16761 294 16780 313
rect 3594 261 3613 280
rect 16563 261 16582 280
rect 16827 261 16846 280
rect 2967 228 2986 247
rect 8346 228 8365 247
rect 13923 228 13942 247
rect 13956 228 13975 247
rect 14319 228 14338 247
rect 14484 228 14503 247
rect 14616 228 14635 247
rect 14913 228 14932 247
rect 15804 228 15823 247
rect 15837 228 15856 247
rect 16134 228 16153 247
rect 16860 228 16879 247
rect 2604 195 2623 214
rect 15408 195 15427 214
rect 15441 195 15460 214
rect 15474 195 15493 214
rect 15507 195 15526 214
rect 15540 195 15559 214
rect 16002 195 16021 214
rect 16596 195 16615 214
rect 16629 195 16648 214
rect 16794 195 16813 214
rect 16827 195 16846 214
rect 16959 195 16978 214
rect 2571 162 2590 181
rect 15738 162 15757 181
rect 16299 162 16318 181
rect 16497 162 16516 181
rect 16530 162 16549 181
rect 2010 129 2029 148
rect 3033 129 3052 148
rect 4056 129 4075 148
rect 7983 129 8002 148
rect 8016 129 8035 148
rect 14286 129 14305 148
rect 15870 129 15889 148
rect 16398 129 16417 148
rect 16431 129 16450 148
rect 16893 129 16912 148
rect 327 96 346 115
rect 1944 96 1963 115
rect 9303 96 9322 115
rect 15936 96 15955 115
rect 15969 96 15988 115
rect 16068 96 16087 115
rect 16101 96 16120 115
rect 16200 96 16219 115
rect 16233 96 16252 115
rect 16365 96 16384 115
rect 16464 96 16483 115
rect 16497 96 16516 115
rect 16827 96 16846 115
rect 16860 96 16879 115
rect 16926 96 16945 115
rect 16959 96 16978 115
rect 16992 96 17011 115
rect 17025 96 17044 115
rect 17124 96 17143 115
rect 13989 63 14008 82
rect 14022 63 14041 82
rect 14979 63 14998 82
rect 15012 63 15031 82
rect 15144 63 15163 82
rect 15177 63 15196 82
rect 17223 63 17242 82
rect 327 30 346 49
rect 13197 30 13216 49
rect 16761 30 16780 49
rect 17124 30 17143 49
rect 294 -3 313 16
rect 13164 -3 13183 16
rect 15375 -3 15394 16
rect 15705 -3 15724 16
rect 16728 -3 16747 16
rect 17091 -3 17110 16
rect 17355 -3 17374 16
rect 294 -960 313 -941
rect 426 -960 445 -941
rect 17157 -960 17176 -941
rect 17289 -960 17308 -941
rect 17421 -960 17440 -941
rect 17553 -960 17572 -941
rect 17619 -960 17638 -941
rect 294 -1686 313 -1667
rect 17190 -993 17209 -974
rect 17322 -993 17341 -974
rect 624 -1026 643 -1007
rect 657 -1026 676 -1007
rect 10986 -1026 11005 -1007
rect 11019 -1026 11038 -1007
rect 17487 -1026 17506 -1007
rect 591 -1059 610 -1040
rect 8940 -1059 8959 -1040
rect 8973 -1059 8992 -1040
rect 657 -1092 676 -1073
rect 690 -1092 709 -1073
rect 822 -1092 841 -1073
rect 855 -1092 874 -1073
rect 12141 -1092 12160 -1073
rect 17322 -1092 17341 -1073
rect 558 -1125 577 -1106
rect 9963 -1125 9982 -1106
rect 9996 -1125 10015 -1106
rect 17190 -1125 17209 -1106
rect 723 -1158 742 -1139
rect 1251 -1158 1270 -1139
rect 1284 -1158 1303 -1139
rect 11019 -1158 11038 -1139
rect 558 -1191 577 -1172
rect 591 -1191 610 -1172
rect 624 -1191 643 -1172
rect 525 -1620 544 -1601
rect 5673 -1191 5692 -1172
rect 5706 -1191 5725 -1172
rect 6696 -1191 6715 -1172
rect 6729 -1191 6748 -1172
rect 9996 -1191 10015 -1172
rect 690 -1224 709 -1205
rect 723 -1224 742 -1205
rect 8973 -1224 8992 -1205
rect 7719 -1257 7738 -1238
rect 6729 -1290 6748 -1271
rect 855 -1323 874 -1304
rect 5706 -1323 5725 -1304
rect 591 -1653 610 -1634
rect 624 -1653 643 -1634
rect 657 -1653 676 -1634
rect 690 -1653 709 -1634
rect 723 -1653 742 -1634
rect 756 -1653 775 -1634
rect 789 -1653 808 -1634
rect 822 -1653 841 -1634
rect 855 -1653 874 -1634
rect 888 -1653 907 -1634
rect 261 -1719 280 -1700
rect 492 -1686 511 -1667
rect 558 -1686 577 -1667
rect 1284 -1356 1303 -1337
rect 360 -1719 379 -1700
rect 657 -1719 676 -1700
rect 888 -1719 907 -1700
rect 294 -1752 313 -1733
rect 327 -1752 346 -1733
rect 261 -1785 280 -1766
rect 855 -1785 874 -1766
rect 327 -1818 346 -1799
rect 360 -1818 379 -1799
rect 393 -1818 412 -1799
rect 822 -1818 841 -1799
rect 426 -1851 445 -1832
rect 459 -1851 478 -1832
rect 789 -1851 808 -1832
rect 294 -1884 313 -1865
rect 327 -1884 346 -1865
rect 360 -1884 379 -1865
rect 756 -1884 775 -1865
rect 261 -1917 280 -1898
rect 723 -1917 742 -1898
rect 690 -1950 709 -1931
rect 162 -1983 181 -1964
rect 195 -1983 214 -1964
rect 228 -1983 247 -1964
<< metal2 >>
rect 330 49 344 96
rect 297 -33 311 -3
rect 1947 -33 1961 96
rect 2013 -33 2027 129
rect 2574 -33 2588 162
rect 2607 -33 2621 195
rect 2970 -33 2984 228
rect 3036 -33 3050 129
rect 3597 -33 3611 261
rect 3630 -33 3644 294
rect 3993 -33 4007 327
rect 4059 -33 4073 129
rect 4620 -33 4634 360
rect 4653 -33 4667 393
rect 5016 -33 5030 426
rect 5082 -33 5096 459
rect 6039 -33 6053 492
rect 6105 -33 6119 525
rect 7062 -33 7076 426
rect 7128 -33 7142 525
rect 7854 -33 7868 558
rect 7887 -33 7901 591
rect 7953 -33 7967 624
rect 8019 148 8033 624
rect 7986 -33 8000 129
rect 8283 -33 8297 624
rect 8349 -33 8363 228
rect 9306 -33 9320 96
rect 9372 -33 9386 657
rect 10329 -33 10343 690
rect 10395 -33 10409 723
rect 11121 -33 11135 756
rect 11220 610 11234 756
rect 11187 -33 11201 591
rect 11484 -33 11498 426
rect 11550 -33 11564 756
rect 12507 -33 12521 789
rect 12573 -33 12587 822
rect 13200 49 13214 822
rect 13167 -33 13181 -3
rect 13299 -33 13313 822
rect 13332 -33 13346 855
rect 13398 -33 13412 888
rect 13464 610 13478 888
rect 13431 -33 13445 591
rect 13497 -33 13511 888
rect 13530 -33 13544 558
rect 13629 478 13643 888
rect 13596 -33 13610 459
rect 13662 -33 13676 888
rect 13794 544 13808 888
rect 13695 -33 13709 459
rect 13761 -33 13775 525
rect 13827 -33 13841 525
rect 13860 -33 13874 888
rect 13959 247 13973 888
rect 14058 643 14072 855
rect 13926 -33 13940 228
rect 14025 82 14039 624
rect 13992 -33 14006 63
rect 14025 -33 14039 63
rect 14091 -33 14105 822
rect 14157 -33 14171 756
rect 14256 478 14270 789
rect 14421 676 14435 756
rect 14223 -33 14237 459
rect 14289 -33 14303 129
rect 14322 -33 14336 228
rect 14388 -33 14402 657
rect 14454 -33 14468 558
rect 14487 -33 14501 228
rect 14553 -33 14567 723
rect 14619 -33 14633 228
rect 14652 -33 14666 492
rect 14718 -33 14732 657
rect 14784 -33 14798 591
rect 14883 478 14897 657
rect 14850 -33 14864 459
rect 14916 -33 14930 228
rect 15015 82 15029 624
rect 14982 -33 14996 63
rect 15048 -33 15062 624
rect 15081 -33 15095 426
rect 15180 82 15194 624
rect 15147 -33 15161 63
rect 15213 -33 15227 624
rect 15345 544 15359 624
rect 15246 -33 15260 459
rect 15312 -33 15326 525
rect 15444 214 15458 591
rect 15510 214 15524 558
rect 15378 -33 15392 -3
rect 15411 -33 15425 195
rect 15477 -33 15491 195
rect 15543 -33 15557 195
rect 15576 -33 15590 492
rect 15675 346 15689 525
rect 15642 -33 15656 327
rect 15840 247 15854 492
rect 15708 -33 15722 -3
rect 15741 -33 15755 162
rect 15807 -33 15821 228
rect 15873 -33 15887 129
rect 15972 115 15986 459
rect 15939 -33 15953 96
rect 16005 -33 16019 195
rect 16104 115 16118 426
rect 16071 -33 16085 96
rect 16137 -33 16151 228
rect 16236 115 16250 393
rect 16203 -33 16217 96
rect 16269 -33 16283 294
rect 16302 -33 16316 162
rect 16434 148 16448 360
rect 16533 181 16547 327
rect 16368 -33 16382 96
rect 16401 -33 16415 129
rect 16500 115 16514 162
rect 16467 -33 16481 96
rect 16500 -33 16514 96
rect 16566 -33 16580 261
rect 16632 214 16646 294
rect 16599 -33 16613 195
rect 16665 -33 16679 294
rect 16764 49 16778 294
rect 16830 214 16844 261
rect 16731 -33 16745 -3
rect 16797 -33 16811 195
rect 16863 115 16877 228
rect 16830 -33 16844 96
rect 16896 -33 16910 129
rect 16962 115 16976 195
rect 16929 -33 16943 96
rect 16995 -33 17009 96
rect 17028 -33 17042 96
rect 17127 49 17141 96
rect 17094 -33 17108 -3
rect 17226 -33 17240 63
rect 17358 -33 17372 -3
rect 297 -941 311 -899
rect 429 -941 443 -899
rect 561 -1172 575 -1125
rect 594 -1172 608 -1059
rect 627 -1172 641 -1026
rect 660 -1073 674 -1026
rect 825 -1073 839 -899
rect 693 -1205 707 -1092
rect 726 -1205 740 -1158
rect 858 -1304 872 -1092
rect 1254 -1139 1268 -899
rect 1287 -1337 1301 -1158
rect 5676 -1172 5690 -899
rect 6699 -1172 6713 -899
rect 5709 -1304 5723 -1191
rect 6732 -1271 6746 -1191
rect 7722 -1238 7736 -899
rect 8943 -1040 8957 -899
rect 8976 -1205 8990 -1059
rect 9966 -1106 9980 -899
rect 10989 -1007 11003 -899
rect 9999 -1172 10013 -1125
rect 11022 -1139 11036 -1026
rect 12144 -1073 12158 -899
rect 17160 -941 17174 -899
rect 17292 -941 17306 -899
rect 17424 -941 17438 -899
rect 17193 -1106 17207 -993
rect 17325 -1073 17339 -993
rect 17490 -1007 17504 -899
rect 17556 -941 17570 -899
rect 17622 -941 17636 -899
rect 264 -1766 278 -1719
rect 297 -1733 311 -1686
rect 330 -1799 344 -1752
rect 363 -1799 377 -1719
rect 165 -2000 179 -1983
rect 198 -2000 212 -1983
rect 231 -2000 245 -1983
rect 264 -2000 278 -1917
rect 297 -2000 311 -1884
rect 330 -2000 344 -1884
rect 363 -2000 377 -1884
rect 396 -2000 410 -1818
rect 429 -2000 443 -1851
rect 462 -2000 476 -1851
rect 495 -2000 509 -1686
rect 528 -2000 542 -1620
rect 561 -2000 575 -1686
rect 594 -2000 608 -1653
rect 627 -2000 641 -1653
rect 660 -1700 674 -1653
rect 693 -1931 707 -1653
rect 726 -1898 740 -1653
rect 759 -1865 773 -1653
rect 792 -1832 806 -1653
rect 825 -1799 839 -1653
rect 858 -1766 872 -1653
rect 891 -1700 905 -1653
use leftbuf  leftbuf_0
timestamp 1673624206
transform 1 0 33 0 1 -899
box 0 0 1650 866
use scanreg  state_reg_2
timestamp 1673624206
transform 1 0 1683 0 1 -899
box 0 0 1023 866
use scanreg  state_reg_0
timestamp 1673624206
transform 1 0 2706 0 1 -899
box 0 0 1023 866
use scanreg  state_reg_1
timestamp 1673624206
transform 1 0 3729 0 1 -899
box 0 0 1023 866
use scanreg  EnableOp1_reg
timestamp 1673624206
transform 1 0 4752 0 1 -899
box 0 0 1023 866
use scanreg  EnableZero_reg
timestamp 1673624206
transform 1 0 5775 0 1 -899
box 0 0 1023 866
use scanreg  LoadA_reg
timestamp 1673624206
transform 1 0 6798 0 1 -899
box 0 0 1023 866
use nand3  g442__2398
timestamp 1673624206
transform 1 0 7821 0 1 -899
box 0 0 198 866
use scanreg  LoadM_reg
timestamp 1673624206
transform 1 0 8019 0 1 -899
box 0 0 1023 866
use scanreg  LoadResult_reg
timestamp 1673624206
transform 1 0 9042 0 1 -899
box 0 0 1023 866
use scanreg  EnableSub_reg
timestamp 1673624206
transform 1 0 10065 0 1 -899
box 0 0 1023 866
use inv  g450
timestamp 1673624206
transform 1 0 11088 0 1 -899
box 0 0 132 866
use scanreg  EnableOp2_reg
timestamp 1673624206
transform 1 0 11220 0 1 -899
box 0 0 1023 866
use scanreg  Done_reg
timestamp 1673624206
transform 1 0 12243 0 1 -899
box 0 0 1023 866
use nand3  g451__5107
timestamp 1673624206
transform 1 0 13266 0 1 -899
box 0 0 198 866
use nand2  g453__6260
timestamp 1673624206
transform 1 0 13464 0 1 -899
box 0 0 165 866
use nand2  g452__4319
timestamp 1673624206
transform 1 0 13629 0 1 -899
box 0 0 165 866
use nand2  g454__8428
timestamp 1673624206
transform 1 0 13794 0 1 -899
box 0 0 165 866
use nand2  g456__5526
timestamp 1673624206
transform 1 0 13959 0 1 -899
box 0 0 165 866
use inv  g458
timestamp 1673624206
transform 1 0 14124 0 1 -899
box 0 0 132 866
use nand2  g460__6783
timestamp 1673624206
transform 1 0 14256 0 1 -899
box 0 0 165 866
use nand2  g461__3680
timestamp 1673624206
transform 1 0 14421 0 1 -899
box 0 0 165 866
use nand2  g462__1617
timestamp 1673624206
transform 1 0 14586 0 1 -899
box 0 0 165 866
use inv  g463
timestamp 1673624206
transform 1 0 14751 0 1 -899
box 0 0 132 866
use inv  g464
timestamp 1673624206
transform 1 0 14883 0 1 -899
box 0 0 132 866
use nand2  g455__2802
timestamp 1673624206
transform 1 0 15015 0 1 -899
box 0 0 165 866
use nand2  g457__1705
timestamp 1673624206
transform 1 0 15180 0 1 -899
box 0 0 165 866
use nand2  g465__5122
timestamp 1673624206
transform 1 0 15345 0 1 -899
box 0 0 165 866
use nand2  g459__8246
timestamp 1673624206
transform 1 0 15510 0 1 -899
box 0 0 165 866
use nand2  g466__7098
timestamp 1673624206
transform 1 0 15675 0 1 -899
box 0 0 165 866
use inv  g467
timestamp 1673624206
transform 1 0 15840 0 1 -899
box 0 0 132 866
use inv  g468
timestamp 1673624206
transform 1 0 15972 0 1 -899
box 0 0 132 866
use inv  g469
timestamp 1673624206
transform 1 0 16104 0 1 -899
box 0 0 132 866
use nand3  g470__6131
timestamp 1673624206
transform 1 0 16236 0 1 -899
box 0 0 198 866
use nand3  g471__1881
timestamp 1673624206
transform 1 0 16434 0 1 -899
box 0 0 198 866
use inv  g473
timestamp 1673624206
transform 1 0 16632 0 1 -899
box 0 0 132 866
use nand3  g472__5115
timestamp 1673624206
transform 1 0 16764 0 1 -899
box 0 0 198 866
use nand2  g474__7482
timestamp 1673624206
transform 1 0 16962 0 1 -899
box 0 0 165 866
use inv  g475
timestamp 1673624206
transform 1 0 17127 0 1 -899
box 0 0 132 866
use inv  g478
timestamp 1673624206
transform 1 0 17259 0 1 -899
box 0 0 132 866
use buffer  rm_assigns_buf_Increment
timestamp 1673624206
transform 1 0 17391 0 1 -899
box 0 0 132 866
use buffer  rm_assigns_buf_LoadB
timestamp 1673624206
transform 1 0 17523 0 1 -899
box 0 0 132 866
use rightend  rightend_0
timestamp 1673624206
transform 1 0 17655 0 1 -899
box 0 0 495 866
<< labels >>
rlabel metal1 0 33 0 45 3 SDO
rlabel metal1 0 66 0 78 3 Req
rlabel metal1 0 99 0 111 3 Done
rlabel metal2 165 -2000 179 -2000 1 SDI
rlabel metal2 198 -2000 212 -2000 1 nReset
rlabel metal2 231 -2000 245 -2000 1 Clock
rlabel metal2 264 -2000 278 -2000 1 Test
rlabel metal2 297 -2000 311 -2000 1 EnableOp2
rlabel metal2 330 -2000 344 -2000 1 EnableZero
rlabel metal2 363 -2000 377 -2000 1 LoadB
rlabel metal2 396 -2000 410 -2000 1 nBorrow
rlabel metal2 429 -2000 443 -2000 1 EnableOp1
rlabel metal2 462 -2000 476 -2000 1 LoadA
rlabel metal2 495 -2000 509 -2000 1 EnableSub
rlabel metal2 528 -2000 542 -2000 1 LoadResult
rlabel metal2 561 -2000 575 -2000 1 Increment
rlabel metal2 594 -2000 608 -2000 1 LoadM
rlabel metal2 627 -2000 641 -2000 1 Overflow
<< end >>
