magic
tech tsmc180
timestamp 1673624206
<< nwell >>
rect 0 429 429 866
<< polysilicon >>
rect 132 805 141 821
rect 198 805 207 823
rect 363 806 372 822
rect 66 716 75 791
rect 132 716 141 756
rect 198 716 207 756
rect 264 716 273 775
rect 66 162 75 667
rect 132 660 141 667
rect 132 162 141 633
rect 198 162 207 667
rect 264 162 273 667
rect 363 195 372 757
rect 66 70 75 135
rect 132 104 141 135
rect 198 104 207 135
rect 264 106 273 135
rect 363 95 372 170
rect 132 65 141 77
rect 198 54 207 77
rect 363 50 372 68
<< ndiffusion >>
rect 54 135 66 162
rect 75 135 132 162
rect 141 135 156 162
rect 177 135 198 162
rect 207 135 264 162
rect 273 135 290 162
rect 116 77 132 104
rect 141 77 155 104
rect 358 68 363 95
rect 372 68 376 95
<< pdiffusion >>
rect 115 756 132 805
rect 141 756 160 805
rect 344 757 363 806
rect 372 757 393 806
rect 46 667 66 716
rect 75 667 93 716
rect 114 667 132 716
rect 141 667 161 716
rect 182 667 198 716
rect 207 667 226 716
rect 247 667 264 716
rect 273 667 290 716
<< pohmic >>
rect 0 31 429 32
rect 0 30 314 31
rect 0 9 160 30
rect 182 9 230 30
rect 252 10 314 30
rect 336 10 429 31
rect 252 9 429 10
rect 0 7 429 9
<< nohmic >>
rect 0 858 429 859
rect 0 837 168 858
rect 191 837 236 858
rect 259 837 300 858
rect 322 837 429 858
rect 0 834 429 837
<< ntransistor >>
rect 66 135 75 162
rect 132 135 141 162
rect 198 135 207 162
rect 264 135 273 162
rect 132 77 141 104
rect 363 68 372 95
<< ptransistor >>
rect 132 756 141 805
rect 363 757 372 806
rect 66 667 75 716
rect 132 667 141 716
rect 198 667 207 716
rect 264 667 273 716
<< polycontact >>
rect 57 791 81 814
rect 192 756 213 805
rect 263 775 286 800
rect 126 633 147 660
rect 355 170 379 195
rect 191 77 212 104
rect 254 81 278 106
rect 61 46 83 70
rect 128 44 153 65
<< ndiffcontact >>
rect 33 135 54 162
rect 156 135 177 162
rect 290 135 311 162
rect 95 77 116 104
rect 155 77 176 104
rect 337 68 358 95
rect 376 68 397 95
<< pdiffcontact >>
rect 94 756 115 805
rect 160 756 181 805
rect 323 757 344 806
rect 393 757 415 806
rect 25 667 46 716
rect 93 667 114 716
rect 161 667 182 716
rect 226 667 247 716
rect 290 667 311 716
<< psubstratetap >>
rect 160 9 182 30
rect 230 9 252 30
rect 314 10 336 31
<< nsubstratetap >>
rect 168 837 191 858
rect 236 837 259 858
rect 300 837 322 858
<< metal1 >>
rect 0 858 429 859
rect 0 837 168 858
rect 191 837 236 858
rect 259 837 300 858
rect 322 837 429 858
rect 0 834 429 837
rect 98 805 110 834
rect 181 756 192 805
rect 31 730 177 742
rect 31 716 43 730
rect 165 716 177 730
rect 230 716 242 834
rect 328 806 340 834
rect 164 652 176 667
rect 295 652 307 667
rect 164 640 307 652
rect 0 434 429 446
rect 0 401 429 413
rect 0 377 429 389
rect 0 353 429 365
rect 0 329 429 341
rect 37 32 49 135
rect 176 77 191 104
rect 99 32 111 77
rect 295 32 307 135
rect 341 32 353 68
rect 0 31 429 32
rect 0 30 314 31
rect 0 9 160 30
rect 182 9 230 30
rect 252 10 314 30
rect 336 10 429 31
rect 252 9 429 10
rect 0 7 429 9
<< m2contact >>
rect 57 791 81 814
rect 263 775 286 800
rect 396 771 415 791
rect 92 682 93 706
rect 93 682 114 706
rect 126 633 147 660
rect 355 170 379 195
rect 154 162 178 163
rect 154 138 156 162
rect 156 138 177 162
rect 177 138 178 162
rect 254 81 278 106
rect 61 46 83 70
rect 128 44 153 65
rect 378 68 397 95
<< metal2 >>
rect 66 814 80 866
rect 95 191 109 682
rect 132 660 146 866
rect 264 800 278 866
rect 396 791 410 866
rect 95 177 355 191
rect 160 163 174 177
rect 396 117 410 771
rect 383 102 410 117
rect 383 95 397 102
rect 66 0 80 46
rect 132 0 146 44
rect 264 0 278 81
rect 383 61 397 68
rect 383 47 410 61
rect 396 0 410 47
<< labels >>
rlabel metal1 0 434 0 446 3 ScanReturn
rlabel metal1 0 401 0 413 3 Scan
rlabel metal1 0 377 0 389 3 Test
rlabel metal1 0 353 0 365 3 Clock
rlabel metal1 0 329 0 341 3 nReset
rlabel metal1 429 434 429 446 3 ScanReturn
rlabel metal1 429 401 429 413 3 Scan
rlabel metal1 429 377 429 389 3 Test
rlabel metal1 429 353 429 365 3 Clock
rlabel metal1 429 329 429 341 3 nReset
rlabel metal1 429 7 429 32 7 GND!
rlabel metal1 0 7 0 32 3 GND!
rlabel metal2 264 0 278 0 1 I0
rlabel metal2 396 0 410 0 1 Y
rlabel metal2 132 0 146 0 1 S
rlabel metal2 66 0 80 0 1 I1
rlabel metal1 0 834 0 859 3 Vdd!
rlabel metal1 429 834 429 859 7 Vdd!
rlabel metal2 264 866 278 866 5 I0
rlabel metal2 396 866 410 866 5 Y
rlabel metal2 132 866 146 866 5 S
rlabel metal2 66 866 80 866 5 I1
<< end >>
