magic
tech tsmc180
timestamp 1672154672
<< nwell >>
rect 0 429 132 866
<< polysilicon >>
rect 58 759 67 794
rect 58 694 67 710
rect 58 651 67 669
rect 50 229 59 585
rect 50 150 59 202
<< ndiffusion >>
rect 47 202 50 229
rect 59 202 71 229
<< pdiffusion >>
rect 55 710 58 759
rect 67 710 70 759
<< pohmic >>
rect 0 7 58 32
rect 83 7 132 32
<< nohmic >>
rect 0 834 52 859
rect 77 834 132 859
<< ntransistor >>
rect 50 202 59 229
<< ptransistor >>
rect 58 710 67 759
<< polycontact >>
rect 43 669 68 694
rect 44 585 69 612
<< ndiffcontact >>
rect 22 202 47 229
rect 71 202 95 229
<< pdiffcontact >>
rect 30 710 55 759
rect 70 710 95 759
<< psubstratetap >>
rect 58 7 83 32
<< nsubstratetap >>
rect 52 834 77 859
<< metal1 >>
rect 0 834 52 859
rect 77 834 132 859
rect 37 759 49 834
rect 81 690 93 710
rect 68 678 93 690
rect 81 608 93 678
rect 69 596 93 608
rect 0 434 132 446
rect 0 401 132 413
rect 0 377 132 389
rect 0 353 132 365
rect 0 329 132 341
rect 28 32 40 202
rect 0 7 58 32
rect 83 7 132 32
<< m2contact >>
rect 44 585 69 612
rect 84 202 95 229
rect 95 202 113 229
<< metal2 >>
rect 99 229 113 866
rect 99 0 113 202
<< labels >>
rlabel metal1 0 7 0 32 3 GND!
rlabel metal1 132 7 132 32 7 GND!
rlabel metal1 0 434 0 446 3 ScanReturn
rlabel metal1 0 401 0 413 3 Scan
rlabel metal1 132 401 132 413 7 Scan
rlabel metal1 0 377 0 389 3 Test
rlabel metal1 132 377 132 389 7 Test
rlabel metal1 0 353 0 365 3 Clock
rlabel metal1 132 353 132 365 7 Clock
rlabel metal1 0 329 0 341 3 nReset
rlabel metal1 132 329 132 341 7 nReset
rlabel metal1 0 834 0 859 3 Vdd!
rlabel metal1 132 434 132 446 7 ScanReturn
rlabel metal1 132 834 132 859 7 Vdd!
rlabel metal2 99 0 113 0 1 Low
rlabel metal2 99 866 113 866 5 Low
<< end >>
