magic
tech tsmc180
timestamp 1672154672
<< nwell >>
rect 0 429 231 866
<< polysilicon >>
rect 34 794 43 805
rect 70 794 79 805
rect 108 794 117 805
rect 147 794 156 805
rect 185 761 194 805
rect 34 731 43 745
rect 70 731 79 745
rect 108 731 117 745
rect 34 668 43 682
rect 70 668 79 682
rect 34 602 43 619
rect 70 602 79 619
rect 108 602 117 682
rect 147 668 156 745
rect 185 731 194 740
rect 147 608 156 619
rect 34 530 43 553
rect 70 530 79 553
rect 108 530 117 553
rect 34 282 43 505
rect 70 282 79 505
rect 108 282 117 505
rect 34 218 43 255
rect 70 218 79 255
rect 34 161 43 191
rect 70 161 79 191
rect 108 161 117 255
rect 147 249 156 587
rect 147 218 156 228
rect 34 95 43 134
rect 70 95 79 134
rect 108 95 117 134
rect 147 95 156 191
rect 185 161 194 682
rect 185 122 194 134
rect 34 57 43 68
rect 70 57 79 68
rect 108 57 117 68
rect 147 57 156 68
rect 185 57 194 101
<< ndiffusion >>
rect 18 276 34 282
rect 31 255 34 276
rect 43 276 70 282
rect 43 255 46 276
rect 67 255 70 276
rect 79 276 108 282
rect 79 255 83 276
rect 104 255 108 276
rect 117 261 120 282
rect 117 255 141 261
rect 10 212 34 218
rect 31 191 34 212
rect 43 191 70 218
rect 79 212 103 218
rect 79 191 82 212
rect 123 212 147 218
rect 144 191 147 212
rect 156 216 180 218
rect 156 191 159 216
rect 10 155 34 161
rect 31 134 34 155
rect 43 134 70 161
rect 79 134 108 161
rect 117 155 141 161
rect 117 134 120 155
rect 161 155 185 161
rect 182 134 185 155
rect 194 160 218 161
rect 194 134 197 160
rect 10 89 34 95
rect 31 68 34 89
rect 43 89 70 95
rect 43 68 46 89
rect 67 68 70 89
rect 79 89 108 95
rect 79 68 82 89
rect 103 68 108 89
rect 117 89 147 95
rect 117 68 120 89
rect 141 68 147 89
rect 156 89 180 95
rect 156 68 159 89
<< pdiffusion >>
rect 31 745 34 794
rect 43 745 46 794
rect 67 745 70 794
rect 79 773 82 794
rect 103 773 108 794
rect 79 745 108 773
rect 117 745 120 794
rect 142 745 147 794
rect 156 773 159 794
rect 156 745 180 773
rect 10 723 34 731
rect 31 682 34 723
rect 43 682 70 731
rect 79 682 108 731
rect 117 729 133 731
rect 117 682 120 729
rect 10 641 34 668
rect 31 619 34 641
rect 43 619 70 668
rect 79 641 95 668
rect 79 619 82 641
rect 161 703 185 731
rect 182 682 185 703
rect 194 720 218 731
rect 194 682 197 720
rect 122 645 147 668
rect 144 623 147 645
rect 122 619 147 623
rect 156 645 180 668
rect 156 620 159 645
rect 156 619 180 620
rect 31 553 34 602
rect 43 581 46 602
rect 67 581 70 602
rect 43 553 70 581
rect 79 575 108 602
rect 79 553 82 575
rect 103 553 108 575
rect 117 575 133 602
rect 117 553 120 575
<< pohmic >>
rect 0 11 7 32
rect 28 11 231 32
rect 0 7 231 11
<< nohmic >>
rect 0 858 231 859
rect 0 837 11 858
rect 32 837 82 858
rect 103 837 231 858
rect 0 834 231 837
<< ntransistor >>
rect 34 255 43 282
rect 70 255 79 282
rect 108 255 117 282
rect 34 191 43 218
rect 70 191 79 218
rect 147 191 156 218
rect 34 134 43 161
rect 70 134 79 161
rect 108 134 117 161
rect 185 134 194 161
rect 34 68 43 95
rect 70 68 79 95
rect 108 68 117 95
rect 147 68 156 95
<< ptransistor >>
rect 34 745 43 794
rect 70 745 79 794
rect 108 745 117 794
rect 147 745 156 794
rect 34 682 43 731
rect 70 682 79 731
rect 108 682 117 731
rect 34 619 43 668
rect 70 619 79 668
rect 185 682 194 731
rect 147 619 156 668
rect 34 553 43 602
rect 70 553 79 602
rect 108 553 117 602
<< polycontact >>
rect 185 740 206 761
rect 147 587 168 608
rect 26 505 47 530
rect 64 505 85 530
rect 99 505 120 530
rect 147 228 168 249
rect 185 101 206 122
<< ndiffcontact >>
rect 10 255 31 276
rect 46 255 67 276
rect 83 255 104 276
rect 120 261 141 282
rect 10 191 31 212
rect 82 191 103 212
rect 123 191 144 212
rect 159 191 180 216
rect 10 134 31 155
rect 120 134 141 155
rect 161 134 182 155
rect 197 134 218 160
rect 10 68 31 89
rect 46 68 67 89
rect 82 68 103 89
rect 120 68 141 89
rect 159 68 180 89
<< pdiffcontact >>
rect 10 745 31 794
rect 46 745 67 794
rect 82 773 103 794
rect 120 745 142 794
rect 159 773 180 794
rect 10 682 31 723
rect 120 682 142 729
rect 10 619 31 641
rect 82 619 103 641
rect 161 682 182 703
rect 197 682 218 720
rect 122 623 144 645
rect 159 620 180 645
rect 10 553 31 602
rect 46 581 67 602
rect 82 553 103 575
rect 120 553 141 575
<< psubstratetap >>
rect 7 11 28 32
<< nsubstratetap >>
rect 11 837 32 858
rect 82 837 103 858
<< metal1 >>
rect 0 858 231 859
rect 0 837 11 858
rect 32 837 82 858
rect 103 837 231 858
rect 0 834 231 837
rect 10 794 22 834
rect 86 794 98 834
rect 67 745 120 757
rect 161 758 173 773
rect 161 746 185 758
rect 10 723 22 745
rect 161 729 173 746
rect 142 717 173 729
rect 161 716 173 717
rect 10 669 22 682
rect 166 669 178 682
rect 10 657 178 669
rect 10 641 22 657
rect 128 645 140 657
rect 31 628 62 640
rect 50 602 62 628
rect 87 599 99 619
rect 87 587 147 599
rect 128 575 140 587
rect 31 554 82 566
rect 0 434 231 446
rect 0 401 231 413
rect 0 377 231 389
rect 0 353 231 365
rect 0 329 231 341
rect 11 288 100 300
rect 11 276 23 288
rect 88 276 100 288
rect 51 208 63 255
rect 123 243 135 261
rect 88 231 147 243
rect 88 212 100 231
rect 31 196 63 208
rect 10 179 22 191
rect 129 179 141 191
rect 10 167 174 179
rect 10 155 22 167
rect 162 155 174 167
rect 10 120 22 134
rect 126 122 138 134
rect 10 108 98 120
rect 126 110 185 122
rect 10 89 22 108
rect 86 89 98 108
rect 159 89 171 110
rect 10 32 22 68
rect 50 56 62 68
rect 124 56 136 68
rect 50 44 136 56
rect 0 11 7 32
rect 28 11 231 32
rect 0 7 231 11
<< m2contact >>
rect 197 690 218 715
rect 159 620 180 645
rect 26 505 47 530
rect 64 505 85 530
rect 99 505 120 530
rect 159 191 180 216
rect 197 134 218 160
<< metal2 >>
rect 33 530 47 866
rect 66 530 80 866
rect 99 530 113 866
rect 165 645 179 866
rect 198 715 212 866
rect 33 0 47 505
rect 66 0 80 505
rect 99 0 113 505
rect 165 216 179 620
rect 165 0 179 191
rect 198 160 212 690
rect 198 0 212 134
<< labels >>
rlabel metal1 0 7 0 32 3 GND!
rlabel metal1 231 7 231 32 7 GND!
rlabel metal1 0 329 0 341 3 nReset
rlabel metal1 231 329 231 341 7 nReset
rlabel metal1 0 353 0 365 3 Clock
rlabel metal1 231 353 231 365 7 Clock
rlabel metal1 0 377 0 389 3 Test
rlabel metal1 231 377 231 389 7 Test
rlabel metal2 66 0 80 0 1 B
rlabel metal2 33 0 47 0 1 A
rlabel metal2 99 0 113 0 1 Cin
rlabel metal2 33 866 47 866 5 A
rlabel metal2 66 866 80 866 5 B
rlabel metal2 99 866 113 866 5 Cin
rlabel metal2 165 0 179 0 1 Cout
rlabel metal2 165 866 179 866 5 Cout
rlabel metal2 198 0 212 0 1 S
rlabel metal2 198 866 212 866 5 S
rlabel metal1 231 401 231 413 7 Scan
rlabel metal1 0 401 0 413 3 Scan
rlabel metal1 231 434 231 446 7 ScanReturn
rlabel metal1 0 434 0 446 3 ScanReturn
rlabel metal1 0 834 0 859 3 Vdd!
rlabel metal1 231 834 231 859 7 Vdd!
<< end >>
