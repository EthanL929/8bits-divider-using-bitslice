magic
tech tsmc180
timestamp 1672154672
<< nwell >>
rect 0 429 297 866
<< polysilicon >>
rect 146 807 155 818
rect 61 733 70 779
rect 61 659 70 708
rect 101 659 110 771
rect 146 659 155 758
rect 190 744 199 782
rect 190 659 199 695
rect 61 574 70 610
rect 101 574 110 610
rect 61 293 70 525
rect 101 293 110 525
rect 146 489 155 610
rect 190 489 199 610
rect 61 193 70 266
rect 101 193 110 266
rect 146 193 155 464
rect 190 193 199 464
rect 61 127 70 166
rect 61 85 70 102
rect 101 85 110 166
rect 146 86 155 166
rect 190 127 199 166
rect 101 55 110 60
rect 190 81 199 100
rect 146 48 155 59
<< ndiffusion >>
rect 58 266 61 293
rect 70 266 73 293
rect 98 266 101 293
rect 110 266 116 293
rect 58 166 61 193
rect 70 166 101 193
rect 110 166 113 193
rect 139 166 146 193
rect 155 166 190 193
rect 199 166 202 193
rect 185 100 190 127
rect 199 100 202 127
rect 143 59 146 86
rect 155 59 159 86
<< pdiffusion >>
rect 143 758 146 807
rect 155 758 159 807
rect 185 695 190 744
rect 199 695 202 744
rect 58 610 61 659
rect 70 610 73 659
rect 98 610 101 659
rect 110 610 118 659
rect 143 610 146 659
rect 155 610 158 659
rect 183 610 190 659
rect 199 610 202 659
rect 33 525 61 574
rect 70 525 101 574
rect 110 525 116 574
<< pohmic >>
rect 0 7 29 32
rect 54 7 208 32
rect 233 7 297 32
<< nohmic >>
rect 0 834 34 859
rect 59 834 202 859
rect 227 834 244 859
rect 269 834 297 859
<< ntransistor >>
rect 61 266 70 293
rect 101 266 110 293
rect 61 166 70 193
rect 101 166 110 193
rect 146 166 155 193
rect 190 166 199 193
rect 190 100 199 127
rect 146 59 155 86
<< ptransistor >>
rect 146 758 155 807
rect 190 695 199 744
rect 61 610 70 659
rect 101 610 110 659
rect 146 610 155 659
rect 190 610 199 659
rect 61 525 70 574
rect 101 525 110 574
<< polycontact >>
rect 88 771 113 796
rect 60 708 85 733
rect 130 464 155 489
rect 177 464 202 489
rect 61 102 86 127
rect 88 60 113 85
<< ndiffcontact >>
rect 33 266 58 293
rect 73 266 98 293
rect 116 266 141 293
rect 33 166 58 193
rect 113 166 139 193
rect 202 166 227 193
rect 160 100 185 127
rect 202 100 227 127
rect 118 59 143 86
rect 159 59 182 86
<< pdiffcontact >>
rect 118 758 143 807
rect 159 758 184 807
rect 160 695 185 744
rect 202 695 227 744
rect 33 610 58 659
rect 73 610 98 659
rect 118 610 143 659
rect 158 610 183 659
rect 202 610 227 659
rect 8 525 33 574
rect 116 525 141 574
<< psubstratetap >>
rect 29 7 54 32
rect 208 7 233 32
<< nsubstratetap >>
rect 34 834 59 859
rect 202 834 227 859
rect 244 834 269 859
<< metal1 >>
rect 0 834 34 859
rect 59 834 202 859
rect 227 834 244 859
rect 269 834 297 859
rect 9 574 21 834
rect 166 807 178 834
rect 113 771 118 796
rect 202 744 227 834
rect 85 712 160 724
rect 249 683 261 834
rect 42 671 137 683
rect 42 659 54 671
rect 124 659 137 671
rect 164 671 261 683
rect 164 659 176 671
rect 81 513 93 610
rect 122 598 135 610
rect 208 598 220 610
rect 122 586 220 598
rect 141 543 226 560
rect 81 501 259 513
rect 0 434 297 446
rect 0 401 297 413
rect 0 377 297 389
rect 0 353 297 365
rect 0 329 297 341
rect 38 305 137 317
rect 38 293 50 305
rect 125 293 137 305
rect 176 267 259 279
rect 38 193 50 266
rect 37 32 49 166
rect 81 152 93 266
rect 176 254 188 267
rect 113 242 188 254
rect 113 193 125 242
rect 151 210 226 222
rect 151 152 163 210
rect 81 140 163 152
rect 215 127 227 166
rect 86 106 160 118
rect 113 60 118 85
rect 164 32 176 59
rect 215 32 227 100
rect 0 7 29 32
rect 54 7 208 32
rect 233 7 297 32
<< m2contact >>
rect 226 540 250 565
rect 259 495 283 520
rect 130 464 155 489
rect 191 464 202 489
rect 202 464 216 489
rect 259 260 283 285
rect 226 205 250 230
<< metal2 >>
rect 132 489 146 866
rect 198 489 212 866
rect 231 565 245 866
rect 132 0 146 464
rect 198 0 212 464
rect 231 230 245 540
rect 264 520 278 866
rect 264 285 278 495
rect 231 0 245 205
rect 264 0 278 260
<< labels >>
rlabel metal1 0 329 0 341 3 nReset
rlabel metal1 0 353 0 365 3 Clock
rlabel metal1 0 377 0 389 3 Test
rlabel metal1 0 434 0 446 3 ScanReturn
rlabel metal1 0 401 0 413 3 Scan
rlabel metal1 0 834 0 859 3 Vdd!
rlabel metal1 0 7 0 32 3 GND!
rlabel metal2 132 0 146 0 1 A
rlabel metal2 132 866 146 866 5 A
rlabel metal2 198 0 212 0 1 B
rlabel metal2 198 866 212 866 5 B
rlabel metal2 231 0 245 0 1 C
rlabel metal2 231 866 245 866 5 C
rlabel metal1 297 834 297 859 7 Vdd!
rlabel metal1 297 434 297 446 7 ScanReturn
rlabel metal1 297 401 297 413 7 Scan
rlabel metal1 297 377 297 389 7 Test
rlabel metal1 297 353 297 365 7 Clock
rlabel metal1 297 329 297 341 7 nReset
rlabel metal1 297 7 297 32 7 GND!
rlabel metal2 264 0 278 0 1 S
rlabel metal2 264 866 278 866 5 S
<< end >>
